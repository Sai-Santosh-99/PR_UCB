module machine1_logic(

   (* buffer_type = "none" *) input [31:0] inform,  
   (* buffer_type = "none" *) input clk,
   (* buffer_type = "none" *) input s_aresetn,
   (* buffer_type = "none" *) input clk_data,
   (* buffer_type = "none" *) output wire [31:0] Q1_t,
   (* buffer_type = "none" *) output wire float_Q1_valid,
   (* buffer_type = "none" *) output wire [31:0] Q2_t,
   (* buffer_type = "none" *) output wire float_Q2_valid
   
   );
   

endmodule
      